module dcache(
    input VA,
    
);


endmodule