module mmu(
    input logic 
    input logic 
);


endmodule