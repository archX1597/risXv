package bpu_pkg;
    import risXv_macro::*;
    `define HIST_LEN 64
    `define BASE_DEPTH
    `define T0_DEPTH
    `define T1_DEPTH
    `define T2_DEPTH
endpackage;