module itlb_ram_line(

);


endmodule