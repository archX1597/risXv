module mmu(
);


endmodule