module dcache(
    input VA,
    input 
);


endmodule