module icache (
        input  logic clk_i,
        input  logic 
        output output_name,
        inout inout_name );
endmodule