module itlb_control (
    
);

endmodule