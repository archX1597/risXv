import mms_pkg::*;

module tlb(
    input [`]
)


endmodule