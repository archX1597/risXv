module dcache(
    input 
);


endmodule