`define DATA_WD 32
`define INST_WD 32