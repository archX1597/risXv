module dcache(
    input 
);	

endmodule
