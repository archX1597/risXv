
module data_ram_bank0;
endmodule

module data_ram_bank1;
endmodule

module data_ram_bank2;
endmodule

module data_ram_bank3;
endmodule